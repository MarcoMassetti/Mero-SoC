VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_2kbyte_1rw_32x512_8
   CLASS BLOCK ;
   SIZE 483.265 BY 325.395 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.54 0.0 116.92 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.38 0.0 122.76 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.22 0.0 128.6 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  134.06 0.0 134.44 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  139.9 0.0 140.28 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  145.74 0.0 146.12 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.58 0.0 151.96 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.42 0.0 157.8 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.26 0.0 163.64 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.1 0.0 169.48 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.94 0.0 175.32 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.78 0.0 181.16 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.62 0.0 187.0 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.46 0.0 192.84 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  198.3 0.0 198.68 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.14 0.0 204.52 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  209.98 0.0 210.36 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  215.82 0.0 216.2 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.66 0.0 222.04 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.5 0.0 227.88 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.34 0.0 233.72 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  239.18 0.0 239.56 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  245.02 0.0 245.4 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.86 0.0 251.24 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  256.7 0.0 257.08 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.54 0.0 262.92 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  268.38 0.0 268.76 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.22 0.0 274.6 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  280.06 0.0 280.44 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  285.9 0.0 286.28 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  291.74 0.0 292.12 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.58 0.0 297.96 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  303.42 0.0 303.8 0.38 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  81.5 0.0 81.88 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.34 0.0 87.72 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 143.185 0.38 143.565 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 151.585 0.38 151.965 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 157.37 0.38 157.75 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 165.87 0.38 166.25 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 171.51 0.38 171.89 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 180.01 0.38 180.39 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 185.185 0.38 185.565 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 193.585 0.38 193.965 ;
      END
   END addr0[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 39.89 0.38 40.27 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 48.39 0.38 48.77 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.635 0.38 41.015 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.18 0.0 93.56 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.02 0.0 99.4 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.86 0.0 105.24 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.7 0.0 111.08 0.38 ;
      END
   END wmask0[3]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  309.26 0.0 309.64 0.38 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.745 0.0 149.125 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  158.49 0.0 158.87 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.295 0.0 167.675 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.49 0.0 178.87 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  188.49 0.0 188.87 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.99 0.0 199.37 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.175 0.0 208.555 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.49 0.0 218.87 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.87 0.0 230.25 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  237.375 0.0 237.755 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.49 0.0 248.87 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  258.49 0.0 258.87 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.07 0.0 269.45 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.255 0.0 278.635 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  288.49 0.0 288.87 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  298.49 0.0 298.87 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  307.225 0.0 307.605 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.49 0.0 318.87 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.49 0.0 328.87 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  338.49 0.0 338.87 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.49 0.0 348.87 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  358.49 0.0 358.87 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  368.49 0.0 368.87 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  378.49 0.0 378.87 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  389.87 0.0 390.25 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  398.49 0.0 398.87 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  408.49 0.0 408.87 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  418.49 0.0 418.87 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  482.885 61.41 483.265 61.79 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  482.885 62.1 483.265 62.48 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  482.885 62.79 483.265 63.17 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  482.885 64.28 483.265 64.66 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  482.885 63.535 483.265 63.915 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 323.655 483.265 325.395 ;
         LAYER met4 ;
         RECT  481.525 0.0 483.265 325.395 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 325.395 ;
         LAYER met3 ;
         RECT  0.0 0.0 483.265 1.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  478.045 3.48 479.785 321.915 ;
         LAYER met3 ;
         RECT  3.48 3.48 479.785 5.22 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 321.915 ;
         LAYER met3 ;
         RECT  3.48 320.175 479.785 321.915 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 482.645 324.775 ;
   LAYER  met2 ;
      RECT  0.62 0.62 482.645 324.775 ;
   LAYER  met3 ;
      RECT  0.98 142.585 482.645 144.165 ;
      RECT  0.62 144.165 0.98 150.985 ;
      RECT  0.62 152.565 0.98 156.77 ;
      RECT  0.62 158.35 0.98 165.27 ;
      RECT  0.62 166.85 0.98 170.91 ;
      RECT  0.62 172.49 0.98 179.41 ;
      RECT  0.62 180.99 0.98 184.585 ;
      RECT  0.62 186.165 0.98 192.985 ;
      RECT  0.62 49.37 0.98 142.585 ;
      RECT  0.62 41.615 0.98 47.79 ;
      RECT  0.98 60.81 482.285 62.39 ;
      RECT  0.98 62.39 482.285 142.585 ;
      RECT  482.285 65.26 482.645 142.585 ;
      RECT  0.62 194.565 0.98 323.055 ;
      RECT  0.62 2.34 0.98 39.29 ;
      RECT  482.285 2.34 482.645 60.81 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 60.81 ;
      RECT  2.88 2.34 480.385 2.88 ;
      RECT  2.88 5.82 480.385 60.81 ;
      RECT  480.385 2.34 482.285 2.88 ;
      RECT  480.385 2.88 482.285 5.82 ;
      RECT  480.385 5.82 482.285 60.81 ;
      RECT  0.98 144.165 2.88 319.575 ;
      RECT  0.98 319.575 2.88 322.515 ;
      RECT  0.98 322.515 2.88 323.055 ;
      RECT  2.88 144.165 480.385 319.575 ;
      RECT  2.88 322.515 480.385 323.055 ;
      RECT  480.385 144.165 482.645 319.575 ;
      RECT  480.385 319.575 482.645 322.515 ;
      RECT  480.385 322.515 482.645 323.055 ;
   LAYER  met4 ;
      RECT  115.94 0.98 117.52 324.775 ;
      RECT  117.52 0.62 121.78 0.98 ;
      RECT  123.36 0.62 127.62 0.98 ;
      RECT  129.2 0.62 133.46 0.98 ;
      RECT  135.04 0.62 139.3 0.98 ;
      RECT  140.88 0.62 145.14 0.98 ;
      RECT  152.56 0.62 156.82 0.98 ;
      RECT  170.08 0.62 174.34 0.98 ;
      RECT  181.76 0.62 186.02 0.98 ;
      RECT  193.44 0.62 197.7 0.98 ;
      RECT  210.96 0.62 215.22 0.98 ;
      RECT  222.64 0.62 226.9 0.98 ;
      RECT  240.16 0.62 244.42 0.98 ;
      RECT  251.84 0.62 256.1 0.98 ;
      RECT  263.52 0.62 267.78 0.98 ;
      RECT  281.04 0.62 285.3 0.98 ;
      RECT  292.72 0.62 296.98 0.98 ;
      RECT  82.48 0.62 86.74 0.98 ;
      RECT  88.32 0.62 92.58 0.98 ;
      RECT  94.16 0.62 98.42 0.98 ;
      RECT  100.0 0.62 104.26 0.98 ;
      RECT  105.84 0.62 110.1 0.98 ;
      RECT  111.68 0.62 115.94 0.98 ;
      RECT  146.72 0.62 148.145 0.98 ;
      RECT  149.725 0.62 150.98 0.98 ;
      RECT  159.47 0.62 162.66 0.98 ;
      RECT  164.24 0.62 166.695 0.98 ;
      RECT  168.275 0.62 168.5 0.98 ;
      RECT  175.92 0.62 177.89 0.98 ;
      RECT  179.47 0.62 180.18 0.98 ;
      RECT  187.6 0.62 187.89 0.98 ;
      RECT  189.47 0.62 191.86 0.98 ;
      RECT  199.97 0.62 203.54 0.98 ;
      RECT  205.12 0.62 207.575 0.98 ;
      RECT  209.155 0.62 209.38 0.98 ;
      RECT  216.8 0.62 217.89 0.98 ;
      RECT  219.47 0.62 221.06 0.98 ;
      RECT  228.48 0.62 229.27 0.98 ;
      RECT  230.85 0.62 232.74 0.98 ;
      RECT  234.32 0.62 236.775 0.98 ;
      RECT  238.355 0.62 238.58 0.98 ;
      RECT  246.0 0.62 247.89 0.98 ;
      RECT  249.47 0.62 250.26 0.98 ;
      RECT  257.68 0.62 257.89 0.98 ;
      RECT  259.47 0.62 261.94 0.98 ;
      RECT  270.05 0.62 273.62 0.98 ;
      RECT  275.2 0.62 277.655 0.98 ;
      RECT  279.235 0.62 279.46 0.98 ;
      RECT  286.88 0.62 287.89 0.98 ;
      RECT  289.47 0.62 291.14 0.98 ;
      RECT  299.47 0.62 302.82 0.98 ;
      RECT  304.4 0.62 306.625 0.98 ;
      RECT  308.205 0.62 308.66 0.98 ;
      RECT  310.24 0.62 317.89 0.98 ;
      RECT  319.47 0.62 327.89 0.98 ;
      RECT  329.47 0.62 337.89 0.98 ;
      RECT  339.47 0.62 347.89 0.98 ;
      RECT  349.47 0.62 357.89 0.98 ;
      RECT  359.47 0.62 367.89 0.98 ;
      RECT  369.47 0.62 377.89 0.98 ;
      RECT  379.47 0.62 389.27 0.98 ;
      RECT  390.85 0.62 397.89 0.98 ;
      RECT  399.47 0.62 407.89 0.98 ;
      RECT  409.47 0.62 417.89 0.98 ;
      RECT  419.47 0.62 480.925 0.98 ;
      RECT  2.34 0.62 80.9 0.98 ;
      RECT  117.52 0.98 477.445 2.88 ;
      RECT  117.52 2.88 477.445 322.515 ;
      RECT  117.52 322.515 477.445 324.775 ;
      RECT  477.445 0.98 480.385 2.88 ;
      RECT  477.445 322.515 480.385 324.775 ;
      RECT  480.385 0.98 480.925 2.88 ;
      RECT  480.385 2.88 480.925 322.515 ;
      RECT  480.385 322.515 480.925 324.775 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 322.515 ;
      RECT  2.34 322.515 2.88 324.775 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 322.515 5.82 324.775 ;
      RECT  5.82 0.98 115.94 2.88 ;
      RECT  5.82 2.88 115.94 322.515 ;
      RECT  5.82 322.515 115.94 324.775 ;
   END
END    sky130_sram_2kbyte_1rw_32x512_8
END    LIBRARY
